module testbench;
  reg clk, reset, writeORread;
  reg [7:0] inbyte;
  reg [31:0] pa;
  reg [255:0] dataBlock;
  wire [7:0] cacheOutput;
  cacheModule uut(clk, reset,pa, writeORread, inbyte, dataBlock, cacheOutput);
  always #5 clk=~clk;
  initial
  begin
    clk=0; reset=1;//writeORread=0;inbyte=7'd9;dataBlock=256'h123456;pa=32'h9876ABC0;
    #20
pa= 32'h1a25;
#20
pa= 32'h1a29;
#20
pa= 32'h5af7;
#20
pa= 32'h5afb;
#20
pa= 32'h5aff;
#20
pa= 32'h5b03;
#20
pa= 32'h5b07;
#20
pa= 32'h5b0b;
#20
pa= 32'h5b0f;
#20
pa= 32'h5b13;
#20
pa= 32'h5b17;
#20
pa= 32'h5b1b;
#20
pa= 32'hdf2;
#20
pa= 32'hdf6;
#20
pa= 32'hdfa;
#20
pa= 32'hdfe;
#20
pa= 32'he02;
#20
pa= 32'h5bc0;
#20
pa= 32'h33e0;
#20
pa= 32'h33e4;
#20
pa= 32'h33e8;
#20
pa= 32'h4664;
#20
pa= 32'h4668;
#20
pa= 32'h466c;
#20
pa= 32'h4670;
#20
pa= 32'h4674;
#20
pa= 32'h4678;
#20
pa= 32'h467c;
#20
pa= 32'h4680;
#20
pa= 32'h4684;
#20
pa= 32'h944;
#20
pa= 32'hbec;
#20
pa= 32'h2b2d;
#20
pa= 32'h2b31;
#20
pa= 32'h2b35;
#20
pa= 32'h7c4c;
#20
pa= 32'h7c50;
#20
pa= 32'h7c54;
#20
pa= 32'h7c58;
#20
pa= 32'h4150;
#20
pa= 32'h1370;
#20
pa= 32'h27b4;
#20
pa= 32'h27b8;
#20
pa= 32'h27bc;
#20
pa= 32'h27c0;
#20
pa= 32'h27c4;
#20
pa= 32'h27c8;
#20
pa= 32'h27cc;
#20
pa= 32'h27d0;
#20
pa= 32'h27d4;
#20
pa= 32'h27d8;
#20
pa= 32'h27dc;
#20
pa= 32'h27e0;
#20
pa= 32'h45f0;
#20
pa= 32'h45f4;
#20
pa= 32'h45f8;
#20
pa= 32'h45fc;
#20
pa= 32'h3c2b;
#20
pa= 32'h3c2f;
#20
pa= 32'h3c33;
#20
pa= 32'h3c37;
#20
pa= 32'h3c3b;
#20
pa= 32'h3c3f;
#20
pa= 32'h3c43;
#20
pa= 32'ha05;
#20
pa= 32'ha09;
#20
pa= 32'ha0d;
#20
pa= 32'ha11;
#20
pa= 32'ha15;
#20
pa= 32'ha19;
#20
pa= 32'h5e87;
#20
pa= 32'h7103;
#20
pa= 32'h7107;
#20
pa= 32'h710b;
#20
pa= 32'h710f;
#20
pa= 32'h7113;
#20
pa= 32'h7117;
#20
pa= 32'h4e8b;
#20
pa= 32'h4e8f;
#20
pa= 32'h4e93;
#20
pa= 32'h4e97;
#20
pa= 32'h4e9b;
#20
pa= 32'h4e9f;
#20
pa= 32'h4ea3;
#20
pa= 32'h4ea7;
#20
pa= 32'h4eab;
#20
pa= 32'h4eaf;
#20
pa= 32'h35b8;
#20
pa= 32'h35bc;
#20
pa= 32'h35c0;
#20
pa= 32'h35c4;
#20
pa= 32'h35c8;
#20
pa= 32'h6d36;
#20
pa= 32'h6d3a;
#20
pa= 32'h6d3e;
#20
pa= 32'h6d42;
#20
pa= 32'h6d46;
#20
pa= 32'h6d4a;
#20
pa= 32'h6d4e;
#20
pa= 32'h6d52;
#20
pa= 32'h6d56;
#20
pa= 32'h6d5a;
#20
pa= 32'h6d5e;
#20
pa= 32'h6d62;
#20
pa= 32'h6d66;
#20
pa= 32'h204b;
#20
pa= 32'h204f;
#20
pa= 32'h2053;
#20
pa= 32'h2057;
#20
pa= 32'h205b;
#20
pa= 32'h205f;
#20
pa= 32'h2063;
#20
pa= 32'h2067;
#20
pa= 32'h206b;
#20
pa= 32'h16be;
#20
pa= 32'h16c2;
#20
pa= 32'h16c6;
#20
pa= 32'h16ca;
#20
pa= 32'h16ce;
#20
pa= 32'h7df3;
#20
pa= 32'h7df7;
#20
pa= 32'h560e;
#20
pa= 32'h5612;
#20
pa= 32'h5702;
#20
pa= 32'h5706;
#20
pa= 32'h570a;
#20
pa= 32'h570e;
#20
pa= 32'h5712;
#20
pa= 32'h5716;
#20
pa= 32'h571a;
#20
pa= 32'h571e;
#20
pa= 32'h5722;
#20
pa= 32'h5726;
#20
pa= 32'h537f;
#20
pa= 32'h5383;
#20
pa= 32'h5387;
#20
pa= 32'h538b;
#20
pa= 32'h538f;
#20
pa= 32'h5393;
#20
pa= 32'h5397;
#20
pa= 32'h7b9a;
#20
pa= 32'h7b9e;
#20
pa= 32'hb50;
#20
pa= 32'hb54;
#20
pa= 32'hb58;
#20
pa= 32'hb5c;
#20
pa= 32'hb60;
#20
pa= 32'hb64;
#20
pa= 32'hb68;
#20
pa= 32'hb6c;
#20
pa= 32'hb70;
#20
pa= 32'h12a2;
#20
pa= 32'h12a6;
#20
pa= 32'h4ba9;
#20
pa= 32'h16d0;
#20
pa= 32'h502f;
#20
pa= 32'h5033;
#20
pa= 32'h5037;
#20
pa= 32'h503b;
#20
pa= 32'h503f;
#20
pa= 32'h5043;
#20
pa= 32'h5047;
#20
pa= 32'h504b;
#20
pa= 32'h504f;
#20
pa= 32'h5053;
#20
pa= 32'h5057;
#20
pa= 32'h23b7;
#20
pa= 32'h23bb;
#20
pa= 32'h40ce;
#20
pa= 32'h40d2;
#20
pa= 32'h40d6;
#20
pa= 32'h40da;
#20
pa= 32'h40de;
#20
pa= 32'h6409;
#20
pa= 32'h640d;
#20
pa= 32'h6411;
#20
pa= 32'h6415;
#20
pa= 32'h41b8;
#20
pa= 32'h41bc;
#20
pa= 32'h41c0;
#20
pa= 32'h3589;
#20
pa= 32'h358d;
#20
pa= 32'h3591;
#20
pa= 32'h3595;
#20
pa= 32'h2364;
#20
pa= 32'h2368;
#20
pa= 32'h236c;
#20
pa= 32'h1b29;
#20
pa= 32'h1b2d;
#20
pa= 32'h5bb1;
#20
pa= 32'h5bb5;
#20
pa= 32'h5bb9;
#20
pa= 32'h5bbd;
#20
pa= 32'h5bc1;
#20
pa= 32'h5bc5;
#20
pa= 32'h5bc9;
#20
pa= 32'h28e3;
#20
pa= 32'h28e7;
#20
pa= 32'h28eb;
#20
pa= 32'h28ef;
#20
pa= 32'h28f3;
#20
pa= 32'h28f7;
#20
pa= 32'h28fb;
#20
pa= 32'h28ff;
#20
pa= 32'h2903;
#20
pa= 32'h787;
#20
pa= 32'h78b;
#20
pa= 32'h78f;
#20
pa= 32'h793;
#20
pa= 32'h797;
#20
pa= 32'h415;
#20
pa= 32'h419;
#20
pa= 32'h41d;
#20
pa= 32'h421;
#20
pa= 32'h425;
#20
pa= 32'h429;
#20
pa= 32'h42d;
#20
pa= 32'h6cd6;
#20
pa= 32'h6cda;
#20
pa= 32'h6cde;
#20
pa= 32'h6ce2;
#20
pa= 32'h61a5;
#20
pa= 32'h61a9;
#20
pa= 32'h61ad;
#20
pa= 32'h61b1;
#20
pa= 32'h61b5;
#20
pa= 32'h170b;
#20
pa= 32'h170f;
#20
pa= 32'h3c28;
#20
pa= 32'h73f6;
#20
pa= 32'h73fa;
#20
pa= 32'h73fe;
#20
pa= 32'h7402;
#20
pa= 32'h7406;
#20
pa= 32'h740a;
#20
pa= 32'h740e;
#20
pa= 32'h7412;
#20
pa= 32'h7416;
#20
pa= 32'h741a;
#20
pa= 32'h741e;
#20
pa= 32'h3839;
#20
pa= 32'h383d;
#20
pa= 32'h1602;
#20
pa= 32'h1606;
#20
pa= 32'h44cb;
#20
pa= 32'h44cf;
#20
pa= 32'h44d3;
#20
pa= 32'h44d7;
#20
pa= 32'h44db;
#20
pa= 32'h44df;
#20
pa= 32'h44e3;
#20
pa= 32'h44e7;
#20
pa= 32'h44eb;
#20
pa= 32'h44ef;
#20
pa= 32'h44f3;
#20
pa= 32'h44f7;
#20
pa= 32'h44fb;
#20
pa= 32'h44ff;
#20
pa= 32'h4503;
#20
pa= 32'h4507;
#20
pa= 32'h450b;
#20
pa= 32'h450f;
#20
pa= 32'h4513;
#20
pa= 32'h4517;
#20
pa= 32'h451b;
#20
pa= 32'h451f;
#20
pa= 32'h4523;
#20
pa= 32'h4527;
#20
pa= 32'h452b;
#20
pa= 32'h452f;
#20
pa= 32'h4533;
#20
pa= 32'h486b;
#20
pa= 32'h486f;
#20
pa= 32'h4873;
#20
pa= 32'h4877;
#20
pa= 32'h487b;
#20
pa= 32'h487f;
#20
pa= 32'h4883;
#20
pa= 32'h6e8d;
#20
pa= 32'h7ad4;
#20
pa= 32'h6075;
#20
pa= 32'h6079;
#20
pa= 32'h607d;
#20
pa= 32'h3966;
#20
pa= 32'h6a1;
#20
pa= 32'h6a5;
#20
pa= 32'h5d72;
#20
pa= 32'h5d76;
#20
pa= 32'h5d7a;
#20
pa= 32'h5d7e;
#20
pa= 32'h5d82;
#20
pa= 32'h77c0;
#20
pa= 32'h77c4;
#20
pa= 32'h77c8;
#20
pa= 32'h77cc;
#20
pa= 32'h77d0;
#20
pa= 32'h77d4;
#20
pa= 32'h6f65;
#20
pa= 32'h6f69;
#20
pa= 32'h27da;
#20
pa= 32'h27de;
#20
pa= 32'h27e2;
#20
pa= 32'h27e6;
#20
pa= 32'h158d;
#20
pa= 32'h1591;
#20
pa= 32'h1595;
#20
pa= 32'h1599;
#20
pa= 32'h7c3f;
#20
pa= 32'h7c43;
#20
pa= 32'h7c47;
#20
pa= 32'h7c4b;
#20
pa= 32'h7c4f;
#20
pa= 32'h7c53;
#20
pa= 32'h7c57;
#20
pa= 32'h8c6;
#20
pa= 32'h8ca;
#20
pa= 32'h8ce;
#20
pa= 32'h8d2;
#20
pa= 32'h8d6;
#20
pa= 32'h8da;
#20
pa= 32'h8de;
#20
pa= 32'h8e2;
#20
pa= 32'h51d2;
#20
pa= 32'h51d6;
#20
pa= 32'h51da;
#20
pa= 32'h16fa;
#20
pa= 32'h16fe;
#20
pa= 32'h1702;
#20
pa= 32'h1706;
#20
pa= 32'h170a;
#20
pa= 32'h170e;
#20
pa= 32'h1712;
#20
pa= 32'h1716;
#20
pa= 32'h171a;
#20
pa= 32'h171e;
#20
pa= 32'h1722;
#20
pa= 32'h1726;
#20
pa= 32'h12f1;
#20
pa= 32'h12f5;
#20
pa= 32'h12f9;
#20
pa= 32'h12fd;
#20
pa= 32'h1301;
#20
pa= 32'h1305;
#20
pa= 32'h1309;
#20
pa= 32'h4e0b;
#20
pa= 32'h4e0f;
#20
pa= 32'h4e13;
#20
pa= 32'h3855;
#20
pa= 32'h8e3;
#20
pa= 32'h15e;
#20
pa= 32'h162;
#20
pa= 32'h166;
#20
pa= 32'h16a;
#20
pa= 32'h16e;
#20
pa= 32'h172;
#20
pa= 32'h176;
#20
pa= 32'h17a;
#20
pa= 32'h17e;
#20
pa= 32'h3f0d;
#20
pa= 32'h3f11;
#20
pa= 32'h3f15;
#20
pa= 32'h3f19;
#20
pa= 32'h3f1d;
#20
pa= 32'h3f21;
#20
pa= 32'h3f25;
#20
pa= 32'h3f29;
#20
pa= 32'h31f5;
#20
pa= 32'h31f9;
#20
pa= 32'h3149;
#20
pa= 32'h314d;
#20
pa= 32'h3151;
#20
pa= 32'h3155;
#20
pa= 32'h3159;
#20
pa= 32'h315d;
#20
pa= 32'h6512;
#20
pa= 32'h6459;
#20
pa= 32'h645d;
#20
pa= 32'h6461;
#20
pa= 32'h6465;
#20
pa= 32'h27a0;
#20
pa= 32'h27a4;
#20
pa= 32'h7b0;
#20
pa= 32'hd8;
#20
pa= 32'hdc;
#20
pa= 32'h3207;
#20
pa= 32'h320b;
#20
pa= 32'h320f;
#20
pa= 32'h3213;
#20
pa= 32'h3f45;
#20
pa= 32'h1e9c;
#20
pa= 32'h1ea0;
#20
pa= 32'ha84;
#20
pa= 32'ha88;
#20
pa= 32'h268e;
#20
pa= 32'h2692;
#20
pa= 32'h2696;
#20
pa= 32'h269a;
#20
pa= 32'h269e;
#20
pa= 32'h26a2;
#20
pa= 32'h26a6;
#20
pa= 32'h5f6d;
#20
pa= 32'h5f71;
#20
pa= 32'h5f75;
#20
pa= 32'h5f79;
#20
pa= 32'h5f7d;
#20
pa= 32'h5f81;
#20
pa= 32'h5f85;
#20
pa= 32'h5f89;
#20
pa= 32'h5f8d;
#20
pa= 32'h5f91;
#20
pa= 32'h255e;
#20
pa= 32'h2562;
#20
pa= 32'h2566;
#20
pa= 32'h256a;
#20
pa= 32'h51fd;
#20
pa= 32'h5201;
#20
pa= 32'h5205;
#20
pa= 32'h5209;
#20
pa= 32'h520d;
#20
pa= 32'h5211;
#20
pa= 32'h5215;
#20
pa= 32'h5219;
#20
pa= 32'h395a;
#20
pa= 32'h395e;
#20
pa= 32'h3962;
#20
pa= 32'h3966;
#20
pa= 32'h396a;
#20
pa= 32'h396e;
#20
pa= 32'h3972;
#20
pa= 32'h260d;
#20
pa= 32'h2611;
#20
pa= 32'h2615;
#20
pa= 32'h2619;
#20
pa= 32'h21e5;
#20
pa= 32'h21e9;
#20
pa= 32'h21ed;
#20
pa= 32'h21f1;
#20
pa= 32'h21f5;
#20
pa= 32'h21f9;
#20
pa= 32'h21fd;
#20
pa= 32'h2201;
#20
pa= 32'h2205;
#20
pa= 32'h75d7;
#20
pa= 32'h5e23;
#20
pa= 32'h5e27;
#20
pa= 32'h5e2b;
#20
pa= 32'h5e2f;
#20
pa= 32'h5e33;
#20
pa= 32'h5e37;
#20
pa= 32'h5e3b;
#20
pa= 32'h5e3f;
#20
pa= 32'h5e43;
#20
pa= 32'h5e47;
#20
pa= 32'h5e4b;
#20
pa= 32'h5e4f;
#20
pa= 32'h5e53;
#20
pa= 32'h5e57;
#20
pa= 32'h5e5b;
#20
pa= 32'h3fd2;
#20
pa= 32'h5902;
#20
pa= 32'h5906;
#20
pa= 32'h590a;
#20
pa= 32'h590e;
#20
pa= 32'h5912;
#20
pa= 32'h5916;
#20
pa= 32'h591a;
#20
pa= 32'h591e;
#20
pa= 32'h5922;
#20
pa= 32'h5926;
#20
pa= 32'h1053;
#20
pa= 32'h1057;
#20
pa= 32'h105b;
#20
pa= 32'h105f;
#20
pa= 32'h4244;
#20
pa= 32'h4248;
#20
pa= 32'h424c;
#20
pa= 32'h4250;
#20
pa= 32'h4254;
#20
pa= 32'h4258;
#20
pa= 32'h4a04;
#20
pa= 32'h2f50;
#20
pa= 32'h2f54;
#20
pa= 32'h2f58;
#20
pa= 32'h2f5c;
#20
pa= 32'h2f60;
#20
pa= 32'h2f64;
#20
pa= 32'h61e6;
#20
pa= 32'h61ea;
#20
pa= 32'h61ee;
#20
pa= 32'h61f2;
#20
pa= 32'h61f6;
#20
pa= 32'h26da;
#20
pa= 32'h884;
#20
pa= 32'h888;
#20
pa= 32'h88c;
#20
pa= 32'h890;
#20
pa= 32'h4683;
#20
pa= 32'h4687;
#20
pa= 32'h41e0;
#20
pa= 32'h41e4;
#20
pa= 32'h41e8;
#20
pa= 32'h41ec;
#20
pa= 32'h41f0;
#20
pa= 32'h41f4;
#20
pa= 32'h41f8;
#20
pa= 32'h41fc;
#20
pa= 32'h4200;
#20
pa= 32'h260c;
#20
pa= 32'h2610;
#20
pa= 32'h2614;
#20
pa= 32'h4688;
#20
pa= 32'h468c;
#20
pa= 32'h4690;
#20
pa= 32'h4694;
#20
pa= 32'h4698;
#20
pa= 32'h469c;
#20
pa= 32'h46a0;
#20
pa= 32'h46a4;
#20
pa= 32'h46a8;
#20
pa= 32'h46ac;
#20
pa= 32'h7c33;
#20
pa= 32'h7c37;
#20
pa= 32'h7c3b;
#20
pa= 32'h7c3f;
#20
pa= 32'h7c43;
#20
pa= 32'h711f;
#20
pa= 32'h7123;
#20
pa= 32'h40b8;
#20
pa= 32'h40bc;
#20
pa= 32'h40c0;
#20
pa= 32'h40c4;
#20
pa= 32'h40c8;
#20
pa= 32'h40cc;
#20
pa= 32'h40d0;
#20
pa= 32'h40d4;
#20
pa= 32'h40d8;
#20
pa= 32'h40dc;
#20
pa= 32'h40e0;
#20
pa= 32'h40e4;
#20
pa= 32'h40e8;
#20
pa= 32'h40ec;
#20
pa= 32'h40f0;
#20
pa= 32'h39e;
#20
pa= 32'h310;
#20
pa= 32'h314;
#20
pa= 32'h318;
#20
pa= 32'h31c;
#20
pa= 32'h320;
#20
pa= 32'h324;
#20
pa= 32'h328;
#20
pa= 32'h32c;
#20
pa= 32'h330;
#20
pa= 32'h334;
#20
pa= 32'h338;
#20
pa= 32'h33c;
#20
pa= 32'h340;
#20
pa= 32'h344;
#20
pa= 32'h348;
#20
pa= 32'h34c;
#20
pa= 32'h26b7;
#20
pa= 32'h26bb;
#20
pa= 32'h26bf;
#20
pa= 32'h4455;
#20
pa= 32'h4459;
#20
pa= 32'h445d;
#20
pa= 32'h2c1b;
#20
pa= 32'h2c1f;
#20
pa= 32'h2c23;
#20
pa= 32'h2c27;
#20
pa= 32'h2c2b;
#20
pa= 32'h2c2f;
#20
pa= 32'h5a64;
#20
pa= 32'h5a68;
#20
pa= 32'h5a6c;
#20
pa= 32'h5a70;
#20
pa= 32'h5a74;
#20
pa= 32'h5a78;
#20
pa= 32'h2978;
#20
pa= 32'h297c;
#20
pa= 32'h2980;
#20
pa= 32'h2984;
#20
pa= 32'h2988;
#20
pa= 32'h298c;
#20
pa= 32'h2990;
#20
pa= 32'h2994;
#20
pa= 32'h2998;
#20
pa= 32'h1070;
#20
pa= 32'h5d1f;
#20
pa= 32'h5d23;
#20
pa= 32'h5d27;
#20
pa= 32'h5d2b;
#20
pa= 32'h1d08;
#20
pa= 32'h6370;
#20
pa= 32'h1520;
#20
pa= 32'h1524;
#20
pa= 32'h344b;
#20
pa= 32'h344f;
#20
pa= 32'h3453;
#20
pa= 32'h3457;
#20
pa= 32'h345b;
#20
pa= 32'hd3e;
#20
pa= 32'hd42;
#20
pa= 32'hd46;
#20
pa= 32'hd4a;
#20
pa= 32'hd4e;
#20
pa= 32'hb84;
#20
pa= 32'hb88;
#20
pa= 32'h485f;
#20
pa= 32'h4863;
#20
pa= 32'h4867;
#20
pa= 32'h486b;
#20
pa= 32'h486f;
#20
pa= 32'h4873;
#20
pa= 32'h4877;
#20
pa= 32'h487b;
#20
pa= 32'h1edd;
#20
pa= 32'h1003;
#20
pa= 32'h1007;
#20
pa= 32'h100b;
#20
pa= 32'h100f;
#20
pa= 32'h1013;
#20
pa= 32'h1017;
#20
pa= 32'h101b;
#20
pa= 32'h499b;
#20
pa= 32'h499f;
#20
pa= 32'h49a3;
#20
pa= 32'h5489;
#20
pa= 32'h548d;
#20
pa= 32'h1ed7;
#20
pa= 32'h2b19;
#20
pa= 32'heba;
#20
pa= 32'hebe;
#20
pa= 32'hec2;
#20
pa= 32'h7187;
#20
pa= 32'h718b;
#20
pa= 32'h718f;
#20
pa= 32'h7193;
#20
pa= 32'h7197;
#20
pa= 32'h719b;
#20
pa= 32'h719f;
#20
pa= 32'h71a3;
#20
pa= 32'h71a7;
#20
pa= 32'h71ab;
#20
pa= 32'h71af;
#20
pa= 32'h3ad0;
#20
pa= 32'h3ad4;
#20
pa= 32'h3ad8;
#20
pa= 32'h3adc;
#20
pa= 32'h3ae0;
#20
pa= 32'h3ae4;
#20
pa= 32'h2824;
#20
pa= 32'h2828;
#20
pa= 32'h282c;
#20
pa= 32'h2830;
#20
pa= 32'h2834;
#20
pa= 32'h388a;
#20
pa= 32'h388e;
#20
pa= 32'h3892;
#20
pa= 32'h3896;
#20
pa= 32'h389a;
#20
pa= 32'hb8f;
#20
pa= 32'hb93;
#20
pa= 32'hb97;
#20
pa= 32'hb9b;
#20
pa= 32'hb9f;
#20
pa= 32'hba3;
#20
pa= 32'hba7;
#20
pa= 32'hbab;
#20
pa= 32'hbaf;
#20
pa= 32'hbb3;
#20
pa= 32'hbb7;
#20
pa= 32'hbbb;
#20
pa= 32'hbbf;
#20
pa= 32'hbc3;
#20
pa= 32'hbc7;
#20
pa= 32'h2869;
#20
pa= 32'h3691;
#20
pa= 32'h3695;
#20
pa= 32'h3699;
#20
pa= 32'h369d;
#20
pa= 32'h36a1;
#20
pa= 32'h36a5;
#20
pa= 32'h36a9;
#20
pa= 32'h36ad;
#20
pa= 32'h36b1;
#20
pa= 32'h36b5;
#20
pa= 32'h7015;
#20
pa= 32'h4cee;
#20
pa= 32'h4cf2;
#20
pa= 32'h4cf6;
#20
pa= 32'h4cfa;
#20
pa= 32'h4cfe;
#20
pa= 32'h4d02;
#20
pa= 32'h4d06;
#20
pa= 32'ha76;
#20
pa= 32'ha7a;
#20
pa= 32'h5bf6;
#20
pa= 32'h5bfa;
#20
pa= 32'h5bfe;
#20
pa= 32'h1706;
#20
pa= 32'h170a;
#20
pa= 32'h170e;
#20
pa= 32'h1712;
#20
pa= 32'h333b;
#20
pa= 32'h333f;
#20
pa= 32'h46d1;
#20
pa= 32'h46d5;
#20
pa= 32'h46d9;
#20
pa= 32'h46dd;
#20
pa= 32'h46e1;
#20
pa= 32'h46e5;
#20
pa= 32'h4b8;
#20
pa= 32'h4bc;
#20
pa= 32'h19de;
#20
pa= 32'h19e2;
#20
pa= 32'h4e3f;
#20
pa= 32'h4e43;
#20
pa= 32'h4e47;
#20
pa= 32'h4e4b;
#20
pa= 32'h4e4f;
#20
pa= 32'h4e53;
#20
pa= 32'h4e57;
#20
pa= 32'h4e5b;
#20
pa= 32'h4e5f;
#20
pa= 32'h4e63;
#20
pa= 32'h4e67;
#20
pa= 32'h4e6b;
#20
pa= 32'h29ad;
#20
pa= 32'h73ae;
#20
pa= 32'h73b2;
#20
pa= 32'h73b6;
#20
pa= 32'h73ba;
#20
pa= 32'h73be;
#20
pa= 32'h73c2;
#20
pa= 32'h58b4;
#20
pa= 32'h7082;
#20
pa= 32'h7086;
#20
pa= 32'h708a;
#20
pa= 32'h708e;
#20
pa= 32'h7092;
#20
pa= 32'h7096;
#20
pa= 32'h709a;
#20
pa= 32'h709e;
#20
pa= 32'h70a2;
#20
pa= 32'h70a6;
#20
pa= 32'h70aa;
#20
pa= 32'h70ae;
#20
pa= 32'h70b2;
#20
pa= 32'h70b6;
#20
pa= 32'h70ba;
#20
pa= 32'h4d30;
#20
pa= 32'h4d34;
#20
pa= 32'h4d38;
#20
pa= 32'h4d3c;
#20
pa= 32'h4d40;
#20
pa= 32'h4d44;
#20
pa= 32'h4d48;
#20
pa= 32'h4d4c;
#20
pa= 32'h4d50;
#20
pa= 32'h4d54;
#20
pa= 32'h4d58;
#20
pa= 32'h4d5c;
#20
pa= 32'h4d60;
#20
pa= 32'h4d64;
#20
pa= 32'h4d68;
#20
pa= 32'h1974;
#20
pa= 32'h1978;
#20
pa= 32'h197c;
#20
pa= 32'h1980;
#20
pa= 32'h1984;
#20
pa= 32'h1988;
#20
pa= 32'h198c;
#20
pa= 32'h515a;
#20
pa= 32'h4eed;
#20
pa= 32'h4ef1;
#20
pa= 32'h2561;
#20
pa= 32'h95;
#20
pa= 32'h3d2c;
#20
pa= 32'h3d30;
#20
pa= 32'h396b;
#20
pa= 32'h1765;
#20
pa= 32'h1769;
#20
pa= 32'h176d;
#20
pa= 32'h1771;
#20
pa= 32'h1775;
#20
pa= 32'h1779;
#20
pa= 32'h177d;
#20
pa= 32'h1781;
#20
pa= 32'h1785;
#20
pa= 32'h1789;
#20
pa= 32'h51a8;
#20
pa= 32'h51ac;
#20
pa= 32'h51b0;
#20
pa= 32'h3bb5;
#20
pa= 32'h56e;
#20
pa= 32'h572;
#20
pa= 32'h576;
#20
pa= 32'h57a;
#20
pa= 32'h57e;
#20
pa= 32'h582;
#20
pa= 32'h586;
#20
pa= 32'h5f3;
#20
pa= 32'h5f7;
#20
pa= 32'h5fb;
#20
pa= 32'h5ff;
#20
pa= 32'h603;
#20
pa= 32'h607;
#20
pa= 32'hdc0;
#20
pa= 32'hdc4;
#20
pa= 32'hdc8;
#20
pa= 32'hdcc;
#20
pa= 32'hdd0;
#20
pa= 32'h72fb;
#20
pa= 32'h72ff;
#20
pa= 32'h7303;
#20
pa= 32'h7307;
#20
pa= 32'h730b;
#20
pa= 32'h730f;
#20
pa= 32'h2f97;
#20
pa= 32'h2f9b;
#20
pa= 32'h2f9f;
#20
pa= 32'h2fa3;
#20
pa= 32'h7d92;
#20
pa= 32'h7d96;
#20
pa= 32'h7d9a;
#20
pa= 32'h7d9e;
#20
pa= 32'h7da2;
#20
pa= 32'h2b2e;
#20
pa= 32'h2b32;
#20
pa= 32'h2b36;
#20
pa= 32'h2b3a;
#20
pa= 32'h13fb;
#20
pa= 32'h13ff;
#20
pa= 32'h1403;
#20
pa= 32'h3940;
#20
pa= 32'h3944;
#20
pa= 32'h3948;
#20
pa= 32'h394c;
#20
pa= 32'h3950;
#20
pa= 32'h3954;
#20
pa= 32'h3958;
#20
pa= 32'h395c;
#20
pa= 32'h3960;
#20
pa= 32'h3964;
#20
pa= 32'h1351;
#20
pa= 32'h1355;
#20
pa= 32'h1359;
#20
pa= 32'h135d;
#20
pa= 32'h1361;
#20
pa= 32'h1365;
#20
pa= 32'h1369;
#20
pa= 32'h136d;
#20
pa= 32'h1371;
#20
pa= 32'h1375;
#20
pa= 32'h1379;
#20
pa= 32'h137d;
#20
pa= 32'h1381;
#20
pa= 32'h567b;
#20
pa= 32'h567f;
#20
pa= 32'h5683;
#20
pa= 32'h5687;
#20
pa= 32'h7842;
#20
pa= 32'h7846;
#20
pa= 32'h3d63;
#20
pa= 32'h3d67;
#20
pa= 32'h3d6b;
#20
pa= 32'h2344;
#20
pa= 32'h2348;
#20
pa= 32'h6a90;
#20
pa= 32'h6a94;
#20
pa= 32'h6a98;
#20
pa= 32'h6a9c;
#20
pa= 32'h6aa0;
#20
pa= 32'h6aa4;
#20
pa= 32'h6aa8;
#20
pa= 32'h6aac;
#20
pa= 32'h502a;
#20
pa= 32'h502e;
#20
pa= 32'h5032;
#20
pa= 32'h6c13;
#20
pa= 32'h6c17;
#20
pa= 32'h6c1b;
#20
pa= 32'h6c1f;
#20
pa= 32'h6c23;
#20
pa= 32'h3393;
#20
pa= 32'h3397;
#20
pa= 32'h339b;
#20
pa= 32'h339f;
#20
pa= 32'hcd2;
#20
pa= 32'hcd6;
#20
pa= 32'h3de1;
#20
pa= 32'h3de5;
#20
pa= 32'h3de9;
#20
pa= 32'h3ded;
#20
pa= 32'h3df1;
#20
pa= 32'h3df5;
#20
pa= 32'h3df9;
#20
pa= 32'h3dfd;
#20
pa= 32'h3e01;
#20
pa= 32'h3e05;
#20
pa= 32'h3e09;
#20
pa= 32'h3e0d;
#20
pa= 32'h3e11;
#20
pa= 32'h3e15;
#20
pa= 32'h2bfc;
#20
pa= 32'h2c00;
#20
pa= 32'h2c04;
#20
pa= 32'h2c08;
#20
pa= 32'h2c0c;
#20
pa= 32'h2c10;
#20
pa= 32'h2c14;
#20
pa= 32'h2c18;
#20
pa= 32'h2c1c;
#20
pa= 32'h2c20;
#20
pa= 32'h2c24;
#20
pa= 32'h2c28;
#20
pa= 32'h2c2c;
#20
pa= 32'h2c30;
#20
pa= 32'h7001;
#20
pa= 32'h7005;
#20
pa= 32'h8fa;
#20
pa= 32'h8fe;
#20
pa= 32'h902;
#20
pa= 32'h906;
#20
pa= 32'h90a;
#20
pa= 32'h90e;
#20
pa= 32'h912;
#20
pa= 32'h916;
#20
pa= 32'h3f03;
#20
pa= 32'h3f07;
#20
pa= 32'h3f0b;
#20
pa= 32'h4ac6;
#20
pa= 32'h4aca;
#20
pa= 32'h4ace;
#20
pa= 32'h4ad2;
#20
pa= 32'h656;
#20
pa= 32'h65a;
#20
pa= 32'h65e;
#20
pa= 32'h662;
#20
pa= 32'h666;
#20
pa= 32'h66a;
#20
pa= 32'h1324;
#20
pa= 32'h1328;
#20
pa= 32'h6437;
#20
pa= 32'h643b;
#20
pa= 32'h643f;
#20
pa= 32'h6443;
#20
pa= 32'h6447;
#20
pa= 32'h644b;
#20
pa= 32'h644f;
#20
pa= 32'h6453;
#20
pa= 32'h6457;
#20
pa= 32'h645b;
#20
pa= 32'h645f;
#20
pa= 32'h3463;
#20
pa= 32'h3467;
#20
pa= 32'h346b;
#20
pa= 32'h346f;
#20
pa= 32'h3473;
#20
pa= 32'h3477;
#20
pa= 32'h2c9b;
#20
pa= 32'h7c55;
#20
pa= 32'h7c59;
#20
pa= 32'h7c5d;
#20
pa= 32'h7c61;
#20
pa= 32'h7c65;
#20
pa= 32'h7c69;
#20
pa= 32'h7c6d;
#20
pa= 32'h7c71;
#20
pa= 32'h7c75;
#20
pa= 32'h7c79;
#20
pa= 32'h7c7d;
#20
pa= 32'h7c81;
#20
pa= 32'h4137;
#20
pa= 32'h413b;
#20
pa= 32'h413f;
#20
pa= 32'h4143;
#20
pa= 32'h4147;
#20
pa= 32'h414b;
#20
pa= 32'h414f;
#20
pa= 32'h4153;
#20
pa= 32'h4157;
#20
pa= 32'h415b;
#20
pa= 32'h415f;
#20
pa= 32'h1249;
#20
pa= 32'h6aba;
#20
pa= 32'h5562;
#20
pa= 32'h5566;
#20
pa= 32'h556a;
#20
pa= 32'h556e;
#20
pa= 32'h655c;
#20
pa= 32'h6560;
#20
pa= 32'h6564;
#20
pa= 32'h6568;
#20
pa= 32'h656c;
#20
pa= 32'h6570;
#20
pa= 32'h5843;
#20
pa= 32'h5847;
#20
pa= 32'h584b;
#20
pa= 32'h584f;
#20
pa= 32'h5853;
#20
pa= 32'h677e;
#20
pa= 32'h6782;
#20
pa= 32'h6786;
#20
pa= 32'h678a;
#20
pa= 32'h678e;
#20
pa= 32'h6792;
#20
pa= 32'h6796;
#20
pa= 32'h679a;
#20
pa= 32'h59d5;
#20
pa= 32'he7c;
#20
pa= 32'h6e65;
#20
pa= 32'h6e69;
#20
pa= 32'h6e6d;
#20
pa= 32'h6e71;
#20
pa= 32'h6e75;
#20
pa= 32'h6e79;
#20
pa= 32'h6e7d;
#20
pa= 32'h6e81;
#20
pa= 32'h6e85;
#20
pa= 32'h6e89;
#20
pa= 32'h6e8d;
#20
pa= 32'h6e91;
#20
pa= 32'h6e95;
#20
pa= 32'h6e99;
#20
pa= 32'h6e9d;
#20
pa= 32'h6ea1;
#20
pa= 32'h6ea5;
#20
pa= 32'h6ea9;
#20
pa= 32'h57ee;
#20
pa= 32'h57f2;
#20
pa= 32'h57f6;
#20
pa= 32'h57fa;
#20
pa= 32'h57fe;
#20
pa= 32'h5802;
#20
pa= 32'h5806;
#20
pa= 32'h580a;
#20
pa= 32'h580e;
#20
pa= 32'h5812;
#20
pa= 32'h7c04;
#20
pa= 32'h7c08;
#20
pa= 32'h7c0c;
#20
pa= 32'h7c10;
#20
pa= 32'h7c14;
#20
pa= 32'h7c18;
#20
pa= 32'h7c1c;
#20
pa= 32'h7c20;
#20
pa= 32'h7c24;
#20
pa= 32'h7c28;
#20
pa= 32'h7c2c;
#20
pa= 32'h7c30;
#20
pa= 32'h7c34;
#20
pa= 32'h7c38;
#20
pa= 32'h7c3c;
#20
pa= 32'h7c40;
#20
pa= 32'h7c44;
#20
pa= 32'h7c48;
#20
pa= 32'h68a5;
#20
pa= 32'h68a9;
#20
pa= 32'h68ad;
#20
pa= 32'h68b1;
#20
pa= 32'h68b5;
#20
pa= 32'h68b9;
#20
pa= 32'h68bd;
#20
pa= 32'h68c1;
#20
pa= 32'h68c5;
#20
pa= 32'h68c9;
#20
pa= 32'h68cd;
#20
pa= 32'h68d1;
#20
pa= 32'h1d59;
#20
pa= 32'h7340;
#20
pa= 32'h7344;
#20
pa= 32'h7348;
#20
pa= 32'h734c;
#20
pa= 32'h7350;
#20
pa= 32'h7354;
#20
pa= 32'h7358;
#20
pa= 32'h735c;
#20
pa= 32'h7360;
#20
pa= 32'h7364;
#20
pa= 32'h7368;
#20
pa= 32'h589c;
#20
pa= 32'h58a0;
#20
pa= 32'h58a4;
#20
pa= 32'h58a8;
#20
pa= 32'h58ac;
#20
pa= 32'h58b0;
#20
pa= 32'h58b4;
#20
pa= 32'h4c13;
#20
pa= 32'h4c17;
#20
pa= 32'h4c1b;
#20
pa= 32'h4c1f;
#20
pa= 32'h4d30;
#20
pa= 32'h4d34;
#20
pa= 32'h4d38;
#20
pa= 32'h4d3c;
#20
pa= 32'h4d40;
#20
pa= 32'h4d44;
#20
pa= 32'h4d48;
#20
pa= 32'h4d4c;
#20
pa= 32'h4d50;
#20
pa= 32'h4d54;
#20
pa= 32'h4d58;
#20
pa= 32'h4d5c;
#20
pa= 32'h4d60;
#20
pa= 32'h4d64;
#20
pa= 32'h4d68;
#20
pa= 32'h84;
#20
pa= 32'h88;
#20
pa= 32'h8c;
#20
pa= 32'h13d1;
#20
pa= 32'h6c11;
#20
pa= 32'h6c15;
#20
pa= 32'h6c19;
#20
pa= 32'h7ed5;
#20
pa= 32'h7ed9;
#20
pa= 32'h7edd;
#20
pa= 32'h7ee1;
#20
pa= 32'h7ee5;
#20
pa= 32'h7ee9;
#20
pa= 32'h598a;
#20
pa= 32'h598e;
#20
pa= 32'h5992;
#20
pa= 32'h590b;
#20
pa= 32'h590f;
#20
pa= 32'h5913;
#20
pa= 32'h4fdd;
#20
pa= 32'h4fe1;
#20
pa= 32'h48e0;
#20
pa= 32'h48e4;
#20
pa= 32'h48e8;
#20
pa= 32'h48ec;
#20
pa= 32'h48f0;
#20
pa= 32'h4dda;
#20
pa= 32'h4dde;
#20
pa= 32'h4de2;
#20
pa= 32'h4de6;
#20
pa= 32'h4dea;
#20
pa= 32'h4dee;
#20
pa= 32'h4df2;
#20
pa= 32'h4df6;
#20
pa= 32'h4ccb;
#20
pa= 32'h4ccf;
#20
pa= 32'h39e7;
#20
pa= 32'h39eb;
#20
pa= 32'h39ef;
#20
pa= 32'h18b3;
#20
pa= 32'h1954;
#20
pa= 32'h1958;
#20
pa= 32'h195c;
#20
pa= 32'h1960;
#20
pa= 32'h1964;
#20
pa= 32'h1968;
#20
pa= 32'h196c;
#20
pa= 32'h222;
#20
pa= 32'h6dc1;
#20
pa= 32'h6dc5;
#20
pa= 32'h6dc9;
#20
pa= 32'h2810;
#20
pa= 32'h3741;
#20
pa= 32'h49f2;
#20
pa= 32'h49f6;
#20
pa= 32'h49fa;
#20
pa= 32'hc4c;
#20
pa= 32'hc50;
#20
pa= 32'hc54;
#20
pa= 32'hc58;
#20
pa= 32'hc5c;
#20
pa= 32'hc60;
#20
pa= 32'hc64;
#20
pa= 32'h2b95;
#20
pa= 32'h2b99;
#20
pa= 32'h2b9d;
#20
pa= 32'h2ba1;
#20
pa= 32'h2ba5;
#20
pa= 32'h2ba9;
#20
pa= 32'h2bad;
#20
pa= 32'h2bb1;
#20
pa= 32'h3039;
#20
pa= 32'h303d;
#20
pa= 32'h3041;
#20
pa= 32'h3045;
#20
pa= 32'h3049;
#20
pa= 32'h304d;
#20
pa= 32'h3051;
#20
pa= 32'h3055;
#20
pa= 32'h32a1;
#20
pa= 32'h32a5;
#20
pa= 32'h32a9;
#20
pa= 32'h32ad;
#20
pa= 32'h32b1;
#20
pa= 32'h32b5;
#20
pa= 32'h32b9;
#20
pa= 32'h32bd;
#20
pa= 32'h32c1;
#20
pa= 32'h32c5;
#20
pa= 32'h32c9;
#20
pa= 32'h32cd;
#20
pa= 32'h32d1;
#20
pa= 32'h32d5;
#20
pa= 32'h32d9;
#20
pa= 32'h32dd;
#20
pa= 32'h32e1;
#20
pa= 32'h32e5;
#20
pa= 32'h32e9;
#20
pa= 32'h32ed;
#20
pa= 32'h32f1;
#20
pa= 32'h32f5;
#20
pa= 32'h32f9;
#20
pa= 32'ha83;
#20
pa= 32'ha87;
#20
pa= 32'h4f9e;
#20
pa= 32'h7f24;
#20
pa= 32'h7f28;
#20
pa= 32'h1dde;
#20
pa= 32'h1de2;
#20
pa= 32'h1de6;
#20
pa= 32'h5b32;
#20
pa= 32'h43e7;
#20
pa= 32'h43eb;
#20
pa= 32'h43ef;
#20
pa= 32'h43f3;
#20
pa= 32'h43f7;
#20
pa= 32'h43fb;
#20
pa= 32'h43ff;
#20
pa= 32'h4403;
#20
pa= 32'h4407;
#20
pa= 32'h440b;
#20
pa= 32'h440f;
#20
pa= 32'h4413;
#20
pa= 32'h4417;
#20
pa= 32'h441b;
#20
pa= 32'h2e51;
#20
pa= 32'h2e55;
#20
pa= 32'h2e59;
#20
pa= 32'h2e5d;
#20
pa= 32'h2e61;
#20
pa= 32'h2e65;
#20
pa= 32'h2e69;
#20
pa= 32'h2e6d;
#20
pa= 32'h74c1;
#20
pa= 32'h74c5;
#20
pa= 32'h74c9;
#20
pa= 32'h74cd;
#20
pa= 32'h74d1;
#20
pa= 32'h3722;
#20
pa= 32'h3726;
#20
pa= 32'h372a;
#20
pa= 32'h372e;
#20
pa= 32'h3732;
$finish;
  end
endmodule